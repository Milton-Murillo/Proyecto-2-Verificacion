// Code your design here
`include "fifo.sv"
`include "Library.sv"
`include "Router_library.sv"
